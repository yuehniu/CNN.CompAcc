/*
 * convolution layer control module
 * parameter:
 *
 * ports:
 *
 * */
module conv_control

endmodule
