/*--------------------------------------------------
 * This module is a ram buffer for every input
 * feature map.
--------------------------------------------------*/
module left_ram


endmodule
