/*--------------------------------------------------
 * This module is top row reg array buffer for
 * storing top row data of input feature map.
--------------------------------------------------*/
module top_row_reg_array


endmodule
